module and_gate (a, b, y);
    input a, b;
    output y;

    or myand(y, a, b);
endmodule
